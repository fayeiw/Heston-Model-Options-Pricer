module ln_lut(
    input clk,
    input en,
    input signed [6:0] x,     
    output signed [31:0] res // Q8.24 format
);

    reg signed [31:0] ln_out;
    assign res = ln_out;

    always@(posedge clk)
    begin
        if (en)
        begin
            case(x)
                10'd1:  ln_out <= -77261934;
                10'd2:  ln_out <= -65632854;
                10'd3:  ln_out <= -58830279;
                10'd4:  ln_out <= -54003774;
                10'd5:  ln_out <= -50260047;
                10'd6:  ln_out <= -47201199;
                10'd7:  ln_out <= -44614980;
                10'd8:  ln_out <= -42374695;
                10'd9:  ln_out <= -40398623;
                10'd10:  ln_out <= -38630967;
                10'd11:  ln_out <= -37031927;
                10'd12:  ln_out <= -35572119;
                10'd13:  ln_out <= -34229225;
                10'd14:  ln_out <= -32985900;
                10'd15:  ln_out <= -31828391;
                10'd16:  ln_out <= -30745615;
                10'd17:  ln_out <= -29728502;
                10'd18:  ln_out <= -28769543;
                10'd19:  ln_out <= -27862446;
                10'd20:  ln_out <= -27001887;
                10'd21:  ln_out <= -26183324;
                10'd22:  ln_out <= -25402848;
                10'd23:  ln_out <= -24657071;
                10'd24:  ln_out <= -23943039;
                10'd25:  ln_out <= -23258159;
                10'd26:  ln_out <= -22600145;
                10'd27:  ln_out <= -21966967;
                10'd28:  ln_out <= -21356820;
                10'd29:  ln_out <= -20768085;
                10'd30:  ln_out <= -20199311;
                10'd31:  ln_out <= -19649189;
                10'd32:  ln_out <= -19116535;
                10'd33:  ln_out <= -18600272;
                10'd34:  ln_out <= -18099422;
                10'd35:  ln_out <= -17613092;
                10'd36:  ln_out <= -17140463;
                10'd37:  ln_out <= -16680785;
                10'd38:  ln_out <= -16233366;
                10'd39:  ln_out <= -15797569;
                10'd40:  ln_out <= -15372807;
                10'd41:  ln_out <= -14958534;
                10'd42:  ln_out <= -14554244;
                10'd43:  ln_out <= -14159468;
                10'd44:  ln_out <= -13773768;
                10'd45:  ln_out <= -13396736;
                10'd46:  ln_out <= -13027991;
                10'd47:  ln_out <= -12667176;
                10'd48:  ln_out <= -12313959;
                10'd49:  ln_out <= -11968025;
                10'd50:  ln_out <= -11629079;
                10'd51:  ln_out <= -11296847;
                10'd52:  ln_out <= -10971065;
                10'd53:  ln_out <= -10651489;
                10'd54:  ln_out <= -10337887;
                10'd55:  ln_out <= -10030040;
                10'd56:  ln_out <= -9727740;
                10'd57:  ln_out <= -9430790;
                10'd58:  ln_out <= -9139005;
                10'd59:  ln_out <= -8852208;
                10'd60:  ln_out <= -8570231;
                10'd61:  ln_out <= -8292916;
                10'd62:  ln_out <= -8020109;
                10'd63:  ln_out <= -7751668;
                10'd64:  ln_out <= -7487455;
                10'd65:  ln_out <= -7227338;
                10'd66:  ln_out <= -6971192;
                10'd67:  ln_out <= -6718898;
                10'd68:  ln_out <= -6470342;
                10'd69:  ln_out <= -6225415;
                10'd70:  ln_out <= -5984012;
                10'd71:  ln_out <= -5746033;
                10'd72:  ln_out <= -5511383;
                10'd73:  ln_out <= -5279970;
                10'd74:  ln_out <= -5051705;
                10'd75:  ln_out <= -4826504;
                10'd76:  ln_out <= -4604286;
                10'd77:  ln_out <= -4384973;
                10'd78:  ln_out <= -4168489;
                10'd79:  ln_out <= -3954764;
                10'd80:  ln_out <= -3743727;
                10'd81:  ln_out <= -3535312;
                10'd82:  ln_out <= -3329454;
                10'd83:  ln_out <= -3126091;
                10'd84:  ln_out <= -2925164;
                10'd85:  ln_out <= -2726615;
                10'd86:  ln_out <= -2530388;
                10'd87:  ln_out <= -2336429;
                10'd88:  ln_out <= -2144688;
                10'd89:  ln_out <= -1955113;
                10'd90:  ln_out <= -1767656;
                10'd91:  ln_out <= -1582270;
                10'd92:  ln_out <= -1398911;
                10'd93:  ln_out <= -1217534;
                10'd94:  ln_out <= -1038097;
                10'd95:  ln_out <= -860558;
                10'd96:  ln_out <= -684879;
                10'd97:  ln_out <= -511020;
                10'd98:  ln_out <= -338945;
                10'd99:  ln_out <= -168616;
                10'd100:  ln_out <= 0;
                default: ln_out <= -32'hFFFFFFFF;
            endcase
        end
    end
endmodule