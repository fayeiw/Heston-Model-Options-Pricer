module sin_lut(
    input clk,
    input en,
    input signed [9:0] x,     
    output signed [31:0] res // Q8.24 format
);

    reg signed [31:0] sin_out;
    assign res = sin_out;

    always@(posedge clk)
    begin
        if (en)
        begin
            case(x)
                10'd1: sin_out <= 167769;
                10'd2: sin_out <= 335521;
                10'd3: sin_out <= 503240;
                10'd4: sin_out <= 670909;
                10'd5: sin_out <= 838511;
                10'd6: sin_out <= 1006029;
                10'd7: sin_out <= 1173446;
                10'd8: sin_out <= 1340746;
                10'd9: sin_out <= 1507911;
                10'd10: sin_out <= 1674926;
                10'd11: sin_out <= 1841774;
                10'd12: sin_out <= 2008437;
                10'd13: sin_out <= 2174900;
                10'd14: sin_out <= 2341144;
                10'd15: sin_out <= 2507155;
                10'd16: sin_out <= 2672915;
                10'd17: sin_out <= 2838408;
                10'd18: sin_out <= 3003617;
                10'd19: sin_out <= 3168526;
                10'd20: sin_out <= 3333118;
                10'd21: sin_out <= 3497376;
                10'd22: sin_out <= 3661285;
                10'd23: sin_out <= 3824828;
                10'd24: sin_out <= 3987988;
                10'd25: sin_out <= 4150749;
                10'd26: sin_out <= 4313095;
                10'd27: sin_out <= 4475010;
                10'd28: sin_out <= 4636478;
                10'd29: sin_out <= 4797482;
                10'd30: sin_out <= 4958006;
                10'd31: sin_out <= 5118034;
                10'd32: sin_out <= 5277551;
                10'd33: sin_out <= 5436539;
                10'd34: sin_out <= 5594984;
                10'd35: sin_out <= 5752870;
                10'd36: sin_out <= 5910180;
                10'd37: sin_out <= 6066900;
                10'd38: sin_out <= 6223012;
                10'd39: sin_out <= 6378503;
                10'd40: sin_out <= 6533355;
                10'd41: sin_out <= 6687554;
                10'd42: sin_out <= 6841085;
                10'd43: sin_out <= 6993931;
                10'd44: sin_out <= 7146078;
                10'd45: sin_out <= 7297510;
                10'd46: sin_out <= 7448213;
                10'd47: sin_out <= 7598171;
                10'd48: sin_out <= 7747368;
                10'd49: sin_out <= 7895792;
                10'd50: sin_out <= 8043425;
                10'd51: sin_out <= 8190255;
                10'd52: sin_out <= 8336265;
                10'd53: sin_out <= 8481442;
                10'd54: sin_out <= 8625770;
                10'd55: sin_out <= 8769236;
                10'd56: sin_out <= 8911825;
                10'd57: sin_out <= 9053523;
                10'd58: sin_out <= 9194315;
                10'd59: sin_out <= 9334189;
                10'd60: sin_out <= 9473128;
                10'd61: sin_out <= 9611121;
                10'd62: sin_out <= 9748152;
                10'd63: sin_out <= 9884208;
                10'd64: sin_out <= 10019276;
                10'd65: sin_out <= 10153343;
                10'd66: sin_out <= 10286393;
                10'd67: sin_out <= 10418416;
                10'd68: sin_out <= 10549396;
                10'd69: sin_out <= 10679321;
                10'd70: sin_out <= 10808179;
                10'd71: sin_out <= 10935955;
                10'd72: sin_out <= 11062639;
                10'd73: sin_out <= 11188215;
                10'd74: sin_out <= 11312673;
                10'd75: sin_out <= 11436000;
                10'd76: sin_out <= 11558183;
                10'd77: sin_out <= 11679211;
                10'd78: sin_out <= 11799070;
                10'd79: sin_out <= 11917750;
                10'd80: sin_out <= 12035238;
                10'd81: sin_out <= 12151522;
                10'd82: sin_out <= 12266591;
                10'd83: sin_out <= 12380434;
                10'd84: sin_out <= 12493038;
                10'd85: sin_out <= 12604393;
                10'd86: sin_out <= 12714488;
                10'd87: sin_out <= 12823311;
                10'd88: sin_out <= 12930852;
                10'd89: sin_out <= 13037100;
                10'd90: sin_out <= 13142044;
                10'd91: sin_out <= 13245674;
                10'd92: sin_out <= 13347980;
                10'd93: sin_out <= 13448950;
                10'd94: sin_out <= 13548576;
                10'd95: sin_out <= 13646847;
                10'd96: sin_out <= 13743753;
                10'd97: sin_out <= 13839285;
                10'd98: sin_out <= 13933433;
                10'd99: sin_out <= 14026188;
                10'd100: sin_out <= 14117540;
                10'd101: sin_out <= 14207480;
                10'd102: sin_out <= 14296000;
                10'd103: sin_out <= 14383090;
                10'd104: sin_out <= 14468741;
                10'd105: sin_out <= 14552946;
                10'd106: sin_out <= 14635696;
                10'd107: sin_out <= 14716982;
                10'd108: sin_out <= 14796796;
                10'd109: sin_out <= 14875131;
                10'd110: sin_out <= 14951978;
                10'd111: sin_out <= 15027330;
                10'd112: sin_out <= 15101179;
                10'd113: sin_out <= 15173518;
                10'd114: sin_out <= 15244340;
                10'd115: sin_out <= 15313637;
                10'd116: sin_out <= 15381403;
                10'd117: sin_out <= 15447631;
                10'd118: sin_out <= 15512314;
                10'd119: sin_out <= 15575446;
                10'd120: sin_out <= 15637021;
                10'd121: sin_out <= 15697031;
                10'd122: sin_out <= 15755472;
                10'd123: sin_out <= 15812338;
                10'd124: sin_out <= 15867622;
                10'd125: sin_out <= 15921319;
                10'd126: sin_out <= 15973425;
                10'd127: sin_out <= 16023933;
                10'd128: sin_out <= 16072839;
                10'd129: sin_out <= 16120137;
                10'd130: sin_out <= 16165823;
                10'd131: sin_out <= 16209893;
                10'd132: sin_out <= 16252342;
                10'd133: sin_out <= 16293166;
                10'd134: sin_out <= 16332360;
                10'd135: sin_out <= 16369921;
                10'd136: sin_out <= 16405845;
                10'd137: sin_out <= 16440129;
                10'd138: sin_out <= 16472768;
                10'd139: sin_out <= 16503761;
                10'd140: sin_out <= 16533102;
                10'd141: sin_out <= 16560791;
                10'd142: sin_out <= 16586824;
                10'd143: sin_out <= 16611198;
                10'd144: sin_out <= 16633910;
                10'd145: sin_out <= 16654960;
                10'd146: sin_out <= 16674344;
                10'd147: sin_out <= 16692060;
                10'd148: sin_out <= 16708108;
                10'd149: sin_out <= 16722484;
                10'd150: sin_out <= 16735188;
                10'd151: sin_out <= 16746219;
                10'd152: sin_out <= 16755575;
                10'd153: sin_out <= 16763256;
                10'd154: sin_out <= 16769260;
                10'd155: sin_out <= 16773588;
                10'd156: sin_out <= 16776238;
                10'd157: sin_out <= 16777210;
                10'd158: sin_out <= 16776505;
                10'd159: sin_out <= 16774122;
                10'd160: sin_out <= 16770062;
                10'd161: sin_out <= 16764324;
                10'd162: sin_out <= 16756911;
                10'd163: sin_out <= 16747821;
                10'd164: sin_out <= 16737057;
                10'd165: sin_out <= 16724619;
                10'd166: sin_out <= 16710509;
                10'd167: sin_out <= 16694728;
                10'd168: sin_out <= 16677277;
                10'd169: sin_out <= 16658159;
                10'd170: sin_out <= 16637374;
                10'd171: sin_out <= 16614926;
                10'd172: sin_out <= 16590817;
                10'd173: sin_out <= 16565048;
                10'd174: sin_out <= 16537623;
                10'd175: sin_out <= 16508544;
                10'd176: sin_out <= 16477815;
                10'd177: sin_out <= 16445437;
                10'd178: sin_out <= 16411415;
                10'd179: sin_out <= 16375752;
                10'd180: sin_out <= 16338452;
                10'd181: sin_out <= 16299517;
                10'd182: sin_out <= 16258953;
                10'd183: sin_out <= 16216762;
                10'd184: sin_out <= 16172950;
                10'd185: sin_out <= 16127521;
                10'd186: sin_out <= 16080479;
                10'd187: sin_out <= 16031829;
                10'd188: sin_out <= 15981576;
                10'd189: sin_out <= 15929725;
                10'd190: sin_out <= 15876280;
                10'd191: sin_out <= 15821249;
                10'd192: sin_out <= 15764635;
                10'd193: sin_out <= 15706444;
                10'd194: sin_out <= 15646683;
                10'd195: sin_out <= 15585357;
                10'd196: sin_out <= 15522473;
                10'd197: sin_out <= 15458037;
                10'd198: sin_out <= 15392054;
                10'd199: sin_out <= 15324533;
                10'd200: sin_out <= 15255479;
                10'd201: sin_out <= 15184899;
                10'd202: sin_out <= 15112801;
                10'd203: sin_out <= 15039192;
                10'd204: sin_out <= 14964079;
                10'd205: sin_out <= 14887470;
                10'd206: sin_out <= 14809371;
                10'd207: sin_out <= 14729792;
                10'd208: sin_out <= 14648740;
                10'd209: sin_out <= 14566223;
                10'd210: sin_out <= 14482249;
                10'd211: sin_out <= 14396828;
                10'd212: sin_out <= 14309966;
                10'd213: sin_out <= 14221674;
                10'd214: sin_out <= 14131959;
                10'd215: sin_out <= 14040831;
                10'd216: sin_out <= 13948299;
                10'd217: sin_out <= 13854373;
                10'd218: sin_out <= 13759061;
                10'd219: sin_out <= 13662373;
                10'd220: sin_out <= 13564318;
                10'd221: sin_out <= 13464908;
                10'd222: sin_out <= 13364150;
                10'd223: sin_out <= 13262057;
                10'd224: sin_out <= 13158637;
                10'd225: sin_out <= 13053902;
                10'd226: sin_out <= 12947861;
                10'd227: sin_out <= 12840525;
                10'd228: sin_out <= 12731905;
                10'd229: sin_out <= 12622012;
                10'd230: sin_out <= 12510857;
                10'd231: sin_out <= 12398451;
                10'd232: sin_out <= 12284805;
                10'd233: sin_out <= 12169930;
                10'd234: sin_out <= 12053839;
                10'd235: sin_out <= 11936542;
                10'd236: sin_out <= 11818051;
                10'd237: sin_out <= 11698379;
                10'd238: sin_out <= 11577537;
                10'd239: sin_out <= 11455537;
                10'd240: sin_out <= 11332391;
                10'd241: sin_out <= 11208112;
                10'd242: sin_out <= 11082713;
                10'd243: sin_out <= 10956205;
                10'd244: sin_out <= 10828602;
                10'd245: sin_out <= 10699916;
                10'd246: sin_out <= 10570159;
                10'd247: sin_out <= 10439346;
                10'd248: sin_out <= 10307489;
                10'd249: sin_out <= 10174601;
                10'd250: sin_out <= 10040696;
                10'd251: sin_out <= 9905787;
                10'd252: sin_out <= 9769887;
                10'd253: sin_out <= 9633010;
                10'd254: sin_out <= 9495169;
                10'd255: sin_out <= 9356380;
                10'd256: sin_out <= 9216654;
                10'd257: sin_out <= 9076007;
                10'd258: sin_out <= 8934453;
                10'd259: sin_out <= 8792005;
                10'd260: sin_out <= 8648677;
                10'd261: sin_out <= 8504485;
                10'd262: sin_out <= 8359443;
                10'd263: sin_out <= 8213564;
                10'd264: sin_out <= 8066864;
                10'd265: sin_out <= 7919358;
                10'd266: sin_out <= 7771059;
                10'd267: sin_out <= 7621984;
                10'd268: sin_out <= 7472146;
                10'd269: sin_out <= 7321561;
                10'd270: sin_out <= 7170244;
                10'd271: sin_out <= 7018210;
                10'd272: sin_out <= 6865474;
                10'd273: sin_out <= 6712052;
                10'd274: sin_out <= 6557958;
                10'd275: sin_out <= 6403208;
                10'd276: sin_out <= 6247819;
                10'd277: sin_out <= 6091804;
                10'd278: sin_out <= 5935180;
                10'd279: sin_out <= 5777963;
                10'd280: sin_out <= 5620168;
                10'd281: sin_out <= 5461811;
                10'd282: sin_out <= 5302908;
                10'd283: sin_out <= 5143474;
                10'd284: sin_out <= 4983526;
                10'd285: sin_out <= 4823080;
                10'd286: sin_out <= 4662152;
                10'd287: sin_out <= 4500757;
                10'd288: sin_out <= 4338912;
                10'd289: sin_out <= 4176634;
                10'd290: sin_out <= 4013937;
                10'd291: sin_out <= 3850839;
                10'd292: sin_out <= 3687357;
                10'd293: sin_out <= 3523505;
                10'd294: sin_out <= 3359301;
                10'd295: sin_out <= 3194761;
                10'd296: sin_out <= 3029902;
                10'd297: sin_out <= 2864740;
                10'd298: sin_out <= 2699291;
                10'd299: sin_out <= 2533572;
                10'd300: sin_out <= 2367600;
                10'd301: sin_out <= 2201392;
                10'd302: sin_out <= 2034963;
                10'd303: sin_out <= 1868330;
                10'd304: sin_out <= 1701511;
                10'd305: sin_out <= 1534522;
                10'd306: sin_out <= 1367379;
                10'd307: sin_out <= 1200099;
                10'd308: sin_out <= 1032700;
                10'd309: sin_out <= 865197;
                10'd310: sin_out <= 697607;
                10'd311: sin_out <= 529948;
                10'd312: sin_out <= 362236;
                10'd313: sin_out <= 194488;
                10'd314: sin_out <= 26720;
                10'd315: sin_out <= -141050;
                10'd316: sin_out <= -308806;
                10'd317: sin_out <= -476532;
                10'd318: sin_out <= -644209;
                10'd319: sin_out <= -811823;
                10'd320: sin_out <= -979355;
                10'd321: sin_out <= -1146789;
                10'd322: sin_out <= -1314109;
                10'd323: sin_out <= -1481297;
                10'd324: sin_out <= -1648337;
                10'd325: sin_out <= -1815213;
                10'd326: sin_out <= -1981906;
                10'd327: sin_out <= -2148402;
                10'd328: sin_out <= -2314683;
                10'd329: sin_out <= -2480732;
                10'd330: sin_out <= -2646533;
                10'd331: sin_out <= -2812070;
                10'd332: sin_out <= -2977325;
                10'd333: sin_out <= -3142283;
                10'd334: sin_out <= -3306926;
                10'd335: sin_out <= -3471239;
                10'd336: sin_out <= -3635204;
                10'd337: sin_out <= -3798806;
                10'd338: sin_out <= -3962028;
                10'd339: sin_out <= -4124854;
                10'd340: sin_out <= -4287268;
                10'd341: sin_out <= -4449253;
                10'd342: sin_out <= -4610792;
                10'd343: sin_out <= -4771871;
                10'd344: sin_out <= -4932473;
                10'd345: sin_out <= -5092581;
                10'd346: sin_out <= -5252180;
                10'd347: sin_out <= -5411254;
                10'd348: sin_out <= -5569787;
                10'd349: sin_out <= -5727762;
                10'd350: sin_out <= -5885165;
                10'd351: sin_out <= -6041980;
                10'd352: sin_out <= -6198190;
                10'd353: sin_out <= -6353781;
                10'd354: sin_out <= -6508736;
                10'd355: sin_out <= -6663040;
                10'd356: sin_out <= -6816678;
                10'd357: sin_out <= -6969634;
                10'd358: sin_out <= -7121894;
                10'd359: sin_out <= -7273441;
                10'd360: sin_out <= -7424261;
                10'd361: sin_out <= -7574338;
                10'd362: sin_out <= -7723658;
                10'd363: sin_out <= -7872205;
                10'd364: sin_out <= -8019966;
                10'd365: sin_out <= -8166924;
                10'd366: sin_out <= -8313066;
                10'd367: sin_out <= -8458376;
                10'd368: sin_out <= -8602841;
                10'd369: sin_out <= -8746445;
                10'd370: sin_out <= -8889175;
                10'd371: sin_out <= -9031016;
                10'd372: sin_out <= -9171953;
                10'd373: sin_out <= -9311974;
                10'd374: sin_out <= -9451063;
                10'd375: sin_out <= -9589207;
                10'd376: sin_out <= -9726392;
                10'd377: sin_out <= -9862605;
                10'd378: sin_out <= -9997831;
                10'd379: sin_out <= -10132058;
                10'd380: sin_out <= -10265271;
                10'd381: sin_out <= -10397458;
                10'd382: sin_out <= -10528606;
                10'd383: sin_out <= -10658700;
                10'd384: sin_out <= -10787728;
                10'd385: sin_out <= -10915678;
                10'd386: sin_out <= -11042536;
                10'd387: sin_out <= -11168290;
                10'd388: sin_out <= -11292927;
                10'd389: sin_out <= -11416435;
                10'd390: sin_out <= -11538801;
                10'd391: sin_out <= -11660013;
                10'd392: sin_out <= -11780059;
                10'd393: sin_out <= -11898928;
                10'd394: sin_out <= -12016606;
                10'd395: sin_out <= -12133083;
                10'd396: sin_out <= -12248346;
                10'd397: sin_out <= -12362385;
                10'd398: sin_out <= -12475187;
                10'd399: sin_out <= -12586742;
                10'd400: sin_out <= -12697038;
                10'd401: sin_out <= -12806065;
                10'd402: sin_out <= -12913811;
                10'd403: sin_out <= -13020265;
                10'd404: sin_out <= -13125418;
                10'd405: sin_out <= -13229258;
                10'd406: sin_out <= -13331775;
                10'd407: sin_out <= -13432959;
                10'd408: sin_out <= -13532800;
                10'd409: sin_out <= -13631287;
                10'd410: sin_out <= -13728411;
                10'd411: sin_out <= -13824163;
                10'd412: sin_out <= -13918532;
                10'd413: sin_out <= -14011509;
                10'd414: sin_out <= -14103085;
                10'd415: sin_out <= -14193251;
                10'd416: sin_out <= -14281997;
                10'd417: sin_out <= -14369315;
                10'd418: sin_out <= -14455197;
                10'd419: sin_out <= -14539633;
                10'd420: sin_out <= -14622614;
                10'd421: sin_out <= -14704134;
                10'd422: sin_out <= -14784183;
                10'd423: sin_out <= -14862754;
                10'd424: sin_out <= -14939839;
                10'd425: sin_out <= -15015429;
                10'd426: sin_out <= -15089518;
                10'd427: sin_out <= -15162098;
                10'd428: sin_out <= -15233162;
                10'd429: sin_out <= -15302703;
                10'd430: sin_out <= -15370713;
                10'd431: sin_out <= -15437187;
                10'd432: sin_out <= -15502116;
                10'd433: sin_out <= -15565496;
                10'd434: sin_out <= -15627318;
                10'd435: sin_out <= -15687579;
                10'd436: sin_out <= -15746270;
                10'd437: sin_out <= -15803387;
                10'd438: sin_out <= -15858923;
                10'd439: sin_out <= -15912874;
                10'd440: sin_out <= -15965233;
                10'd441: sin_out <= -16015996;
                10'd442: sin_out <= -16065157;
                10'd443: sin_out <= -16112712;
                10'd444: sin_out <= -16158655;
                10'd445: sin_out <= -16202983;
                10'd446: sin_out <= -16245690;
                10'd447: sin_out <= -16286773;
                10'd448: sin_out <= -16326227;
                10'd449: sin_out <= -16364048;
                10'd450: sin_out <= -16400233;
                10'd451: sin_out <= -16434779;
                10'd452: sin_out <= -16467680;
                10'd453: sin_out <= -16498935;
                10'd454: sin_out <= -16528540;
                10'd455: sin_out <= -16556492;
                10'd456: sin_out <= -16582789;
                10'd457: sin_out <= -16607427;
                10'd458: sin_out <= -16630404;
                10'd459: sin_out <= -16651719;
                10'd460: sin_out <= -16671368;
                10'd461: sin_out <= -16689350;
                10'd462: sin_out <= -16705664;
                10'd463: sin_out <= -16720306;
                10'd464: sin_out <= -16733277;
                10'd465: sin_out <= -16744574;
                10'd466: sin_out <= -16754197;
                10'd467: sin_out <= -16762145;
                10'd468: sin_out <= -16768416;
                10'd469: sin_out <= -16773011;
                10'd470: sin_out <= -16775928;
                10'd471: sin_out <= -16777168;
                10'd472: sin_out <= -16776730;
                10'd473: sin_out <= -16774614;
                10'd474: sin_out <= -16770821;
                10'd475: sin_out <= -16765350;
                10'd476: sin_out <= -16758204;
                10'd477: sin_out <= -16749381;
                10'd478: sin_out <= -16738884;
                10'd479: sin_out <= -16726712;
                10'd480: sin_out <= -16712868;
                10'd481: sin_out <= -16697353;
                10'd482: sin_out <= -16680168;
                10'd483: sin_out <= -16661315;
                10'd484: sin_out <= -16640796;
                10'd485: sin_out <= -16618613;
                10'd486: sin_out <= -16594768;
                10'd487: sin_out <= -16569263;
                10'd488: sin_out <= -16542102;
                10'd489: sin_out <= -16513286;
                10'd490: sin_out <= -16482819;
                10'd491: sin_out <= -16450704;
                10'd492: sin_out <= -16416944;
                10'd493: sin_out <= -16381542;
                10'd494: sin_out <= -16344502;
                10'd495: sin_out <= -16305827;
                10'd496: sin_out <= -16265522;
                10'd497: sin_out <= -16223591;
                10'd498: sin_out <= -16180037;
                10'd499: sin_out <= -16134865;
                10'd500: sin_out <= -16088079;
                10'd501: sin_out <= -16039685;
                10'd502: sin_out <= -15989687;
                10'd503: sin_out <= -15938090;
                10'd504: sin_out <= -15884899;
                10'd505: sin_out <= -15830119;
                10'd506: sin_out <= -15773757;
                10'd507: sin_out <= -15715817;
                10'd508: sin_out <= -15656306;
                10'd509: sin_out <= -15595229;
                10'd510: sin_out <= -15532592;
                10'd511: sin_out <= -15468403;
                10'd512: sin_out <= -15402666;
                10'd513: sin_out <= -15335389;
                10'd514: sin_out <= -15266579;
                10'd515: sin_out <= -15196242;
                10'd516: sin_out <= -15124386;
                10'd517: sin_out <= -15051017;
                10'd518: sin_out <= -14976142;
                10'd519: sin_out <= -14899771;
                10'd520: sin_out <= -14821909;
                10'd521: sin_out <= -14742565;
                10'd522: sin_out <= -14661747;
                10'd523: sin_out <= -14579463;
                10'd524: sin_out <= -14495721;
                10'd525: sin_out <= -14410529;
                10'd526: sin_out <= -14323896;
                10'd527: sin_out <= -14235831;
                10'd528: sin_out <= -14146342;
                10'd529: sin_out <= -14055439;
                10'd530: sin_out <= -13963130;
                10'd531: sin_out <= -13869425;
                10'd532: sin_out <= -13774333;
                10'd533: sin_out <= -13677863;
                10'd534: sin_out <= -13580026;
                10'd535: sin_out <= -13480831;
                10'd536: sin_out <= -13380287;
                10'd537: sin_out <= -13278406;
                10'd538: sin_out <= -13175197;
                10'd539: sin_out <= -13070670;
                10'd540: sin_out <= -12964836;
                10'd541: sin_out <= -12857706;
                10'd542: sin_out <= -12749290;
                10'd543: sin_out <= -12639599;
                10'd544: sin_out <= -12528644;
                10'd545: sin_out <= -12416436;
                10'd546: sin_out <= -12302987;
                10'd547: sin_out <= -12188307;
                10'd548: sin_out <= -12072409;
                10'd549: sin_out <= -11955303;
                10'd550: sin_out <= -11837002;
                10'd551: sin_out <= -11717517;
                10'd552: sin_out <= -11596860;
                10'd553: sin_out <= -11475044;
                10'd554: sin_out <= -11352080;
                10'd555: sin_out <= -11227981;
                10'd556: sin_out <= -11102759;
                10'd557: sin_out <= -10976427;
                10'd558: sin_out <= -10848998;
                10'd559: sin_out <= -10720483;
                10'd560: sin_out <= -10590896;
                10'd561: sin_out <= -10460251;
                10'd562: sin_out <= -10328559;
                10'd563: sin_out <= -10195834;
                10'd564: sin_out <= -10062090;
                10'd565: sin_out <= -9927340;
                10'd566: sin_out <= -9791597;
                10'd567: sin_out <= -9654874;
                10'd568: sin_out <= -9517187;
                10'd569: sin_out <= -9378547;
                10'd570: sin_out <= -9238970;
                10'd571: sin_out <= -9098469;
                10'd572: sin_out <= -8957058;
                10'd573: sin_out <= -8814751;
                10'd574: sin_out <= -8671563;
                10'd575: sin_out <= -8527507;
                10'd576: sin_out <= -8382599;
                10'd577: sin_out <= -8236853;
                10'd578: sin_out <= -8090283;
                10'd579: sin_out <= -7942904;
                10'd580: sin_out <= -7794731;
                10'd581: sin_out <= -7645778;
                10'd582: sin_out <= -7496060;
                10'd583: sin_out <= -7345594;
                10'd584: sin_out <= -7194392;
                10'd585: sin_out <= -7042471;
                10'd586: sin_out <= -6889846;
                10'd587: sin_out <= -6736532;
                10'd588: sin_out <= -6582544;
                10'd589: sin_out <= -6427898;
                10'd590: sin_out <= -6272609;
                10'd591: sin_out <= -6116693;
                10'd592: sin_out <= -5960165;
                10'd593: sin_out <= -5803041;
                10'd594: sin_out <= -5645337;
                10'd595: sin_out <= -5487069;
                10'd596: sin_out <= -5328251;
                10'd597: sin_out <= -5168901;
                10'd598: sin_out <= -5009034;
                10'd599: sin_out <= -4848666;
                10'd600: sin_out <= -4687814;
                10'd601: sin_out <= -4526492;
                10'd602: sin_out <= -4364718;
                10'd603: sin_out <= -4202507;
                10'd604: sin_out <= -4039876;
                10'd605: sin_out <= -3876841;
                10'd606: sin_out <= -3713419;
                10'd607: sin_out <= -3549625;
                10'd608: sin_out <= -3385476;
                10'd609: sin_out <= -3220989;
                10'd610: sin_out <= -3056179;
                10'd611: sin_out <= -2891064;
                10'd612: sin_out <= -2725660;
                10'd613: sin_out <= -2559983;
                10'd614: sin_out <= -2394050;
                10'd615: sin_out <= -2227878;
                10'd616: sin_out <= -2061483;
                10'd617: sin_out <= -1894882;
                10'd618: sin_out <= -1728091;
                10'd619: sin_out <= -1561128;
                10'd620: sin_out <= -1394008;
                10'd621: sin_out <= -1226749;
                10'd622: sin_out <= -1059368;
                10'd623: sin_out <= -891880;
                10'd624: sin_out <= -724304;
                10'd625: sin_out <= -556654;
                10'd626: sin_out <= -388950;
                10'd627: sin_out <= -221206;
                10'd628: sin_out <= -53440;
                default: sin_out <= -32'hFFFFFFFF;
            endcase
        end
    end
endmodule