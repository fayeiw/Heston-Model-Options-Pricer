module sqrt_lut(
    input clk,
    input en,
    input signed [9:0] x,     
    output signed [31:0] res // Q8.24 format
);

    reg signed [31:0] sqrt_out;
    assign res = sqrt_out;

    always@(posedge clk)
    begin
        if (en)
        begin
            case(x)
                10'd1: sqrt_out <= 1677721;
                10'd2: sqrt_out <= 2372656;
                10'd3: sqrt_out <= 2905899;
                10'd4: sqrt_out <= 3355443;
                10'd5: sqrt_out <= 3751499;
                10'd6: sqrt_out <= 4109561;
                10'd7: sqrt_out <= 4438834;
                10'd8: sqrt_out <= 4745313;
                10'd9: sqrt_out <= 5033164;
                10'd10: sqrt_out <= 5305421;
                10'd11: sqrt_out <= 5564373;
                10'd12: sqrt_out <= 5811798;
                10'd13: sqrt_out <= 6049111;
                10'd14: sqrt_out <= 6277459;
                10'd15: sqrt_out <= 6497787;
                10'd16: sqrt_out <= 6710886;
                10'd17: sqrt_out <= 6917423;
                10'd18: sqrt_out <= 7117969;
                10'd19: sqrt_out <= 7313018;
                10'd20: sqrt_out <= 7502999;
                10'd21: sqrt_out <= 7688286;
                10'd22: sqrt_out <= 7869211;
                10'd23: sqrt_out <= 8046070;
                10'd24: sqrt_out <= 8219123;
                10'd25: sqrt_out <= 8388608;
                10'd26: sqrt_out <= 8554735;
                10'd27: sqrt_out <= 8717697;
                10'd28: sqrt_out <= 8877668;
                10'd29: sqrt_out <= 9034807;
                10'd30: sqrt_out <= 9189259;
                10'd31: sqrt_out <= 9341158;
                10'd32: sqrt_out <= 9490626;
                10'd33: sqrt_out <= 9637776;
                10'd34: sqrt_out <= 9782713;
                10'd35: sqrt_out <= 9925534;
                10'd36: sqrt_out <= 10066329;
                10'd37: sqrt_out <= 10205182;
                10'd38: sqrt_out <= 10342170;
                10'd39: sqrt_out <= 10477368;
                10'd40: sqrt_out <= 10610843;
                10'd41: sqrt_out <= 10742659;
                10'd42: sqrt_out <= 10872878;
                10'd43: sqrt_out <= 11001556;
                10'd44: sqrt_out <= 11128746;
                10'd45: sqrt_out <= 11254498;
                10'd46: sqrt_out <= 11378861;
                10'd47: sqrt_out <= 11501879;
                10'd48: sqrt_out <= 11623596;
                10'd49: sqrt_out <= 11744051;
                10'd50: sqrt_out <= 11863283;
                10'd51: sqrt_out <= 11981328;
                10'd52: sqrt_out <= 12098222;
                10'd53: sqrt_out <= 12213997;
                10'd54: sqrt_out <= 12328685;
                10'd55: sqrt_out <= 12442316;
                10'd56: sqrt_out <= 12554918;
                10'd57: sqrt_out <= 12666520;
                10'd58: sqrt_out <= 12777147;
                10'd59: sqrt_out <= 12886824;
                10'd60: sqrt_out <= 12995575;
                10'd61: sqrt_out <= 13103424;
                10'd62: sqrt_out <= 13210393;
                10'd63: sqrt_out <= 13316502;
                10'd64: sqrt_out <= 13421772;
                10'd65: sqrt_out <= 13526223;
                10'd66: sqrt_out <= 13629874;
                10'd67: sqrt_out <= 13732743;
                10'd68: sqrt_out <= 13834846;
                10'd69: sqrt_out <= 13936202;
                10'd70: sqrt_out <= 14036825;
                10'd71: sqrt_out <= 14136733;
                10'd72: sqrt_out <= 14235939;
                10'd73: sqrt_out <= 14334459;
                10'd74: sqrt_out <= 14432306;
                10'd75: sqrt_out <= 14529495;
                10'd76: sqrt_out <= 14626037;
                10'd77: sqrt_out <= 14721947;
                10'd78: sqrt_out <= 14817235;
                10'd79: sqrt_out <= 14911915;
                10'd80: sqrt_out <= 15005998;
                10'd81: sqrt_out <= 15099494;
                10'd82: sqrt_out <= 15192415;
                10'd83: sqrt_out <= 15284771;
                10'd84: sqrt_out <= 15376572;
                10'd85: sqrt_out <= 15467828;
                10'd86: sqrt_out <= 15558550;
                10'd87: sqrt_out <= 15648745;
                10'd88: sqrt_out <= 15738423;
                10'd89: sqrt_out <= 15827593;
                10'd90: sqrt_out <= 15916264;
                10'd91: sqrt_out <= 16004444;
                10'd92: sqrt_out <= 16092140;
                10'd93: sqrt_out <= 16179361;
                10'd94: sqrt_out <= 16266114;
                10'd95: sqrt_out <= 16352407;
                10'd96: sqrt_out <= 16438247;
                10'd97: sqrt_out <= 16523641;
                10'd98: sqrt_out <= 16608596;
                10'd99: sqrt_out <= 16693119;
                10'd100: sqrt_out <= 16777216;
                10'd101: sqrt_out <= 16860893;
                10'd102: sqrt_out <= 16944157;
                10'd103: sqrt_out <= 17027014;
                10'd104: sqrt_out <= 17109470;
                10'd105: sqrt_out <= 17191530;
                10'd106: sqrt_out <= 17273201;
                10'd107: sqrt_out <= 17354487;
                10'd108: sqrt_out <= 17435394;
                10'd109: sqrt_out <= 17515927;
                10'd110: sqrt_out <= 17596092;
                10'd111: sqrt_out <= 17675893;
                10'd112: sqrt_out <= 17755336;
                10'd113: sqrt_out <= 17834425;
                10'd114: sqrt_out <= 17913164;
                10'd115: sqrt_out <= 17991559;
                10'd116: sqrt_out <= 18069614;
                10'd117: sqrt_out <= 18147333;
                10'd118: sqrt_out <= 18224721;
                10'd119: sqrt_out <= 18301781;
                10'd120: sqrt_out <= 18378519;
                10'd121: sqrt_out <= 18454937;
                10'd122: sqrt_out <= 18531040;
                10'd123: sqrt_out <= 18606832;
                10'd124: sqrt_out <= 18682317;
                10'd125: sqrt_out <= 18757497;
                10'd126: sqrt_out <= 18832378;
                10'd127: sqrt_out <= 18906962;
                10'd128: sqrt_out <= 18981253;
                10'd129: sqrt_out <= 19055254;
                10'd130: sqrt_out <= 19128969;
                10'd131: sqrt_out <= 19202401;
                10'd132: sqrt_out <= 19275553;
                10'd133: sqrt_out <= 19348429;
                10'd134: sqrt_out <= 19421031;
                10'd135: sqrt_out <= 19493363;
                10'd136: sqrt_out <= 19565427;
                10'd137: sqrt_out <= 19637227;
                10'd138: sqrt_out <= 19708766;
                10'd139: sqrt_out <= 19780045;
                10'd140: sqrt_out <= 19851069;
                10'd141: sqrt_out <= 19921840;
                10'd142: sqrt_out <= 19992360;
                10'd143: sqrt_out <= 20062632;
                10'd144: sqrt_out <= 20132659;
                10'd145: sqrt_out <= 20202443;
                10'd146: sqrt_out <= 20271987;
                10'd147: sqrt_out <= 20341293;
                10'd148: sqrt_out <= 20410364;
                10'd149: sqrt_out <= 20479202;
                10'd150: sqrt_out <= 20547809;
                10'd151: sqrt_out <= 20616188;
                10'd152: sqrt_out <= 20684341;
                10'd153: sqrt_out <= 20752270;
                10'd154: sqrt_out <= 20819977;
                10'd155: sqrt_out <= 20887465;
                10'd156: sqrt_out <= 20954736;
                10'd157: sqrt_out <= 21021791;
                10'd158: sqrt_out <= 21088633;
                10'd159: sqrt_out <= 21155264;
                10'd160: sqrt_out <= 21221686;
                10'd161: sqrt_out <= 21287900;
                10'd162: sqrt_out <= 21353909;
                10'd163: sqrt_out <= 21419715;
                10'd164: sqrt_out <= 21485319;
                10'd165: sqrt_out <= 21550724;
                10'd166: sqrt_out <= 21615930;
                10'd167: sqrt_out <= 21680941;
                10'd168: sqrt_out <= 21745757;
                10'd169: sqrt_out <= 21810380;
                10'd170: sqrt_out <= 21874813;
                10'd171: sqrt_out <= 21939056;
                10'd172: sqrt_out <= 22003112;
                10'd173: sqrt_out <= 22066982;
                10'd174: sqrt_out <= 22130667;
                10'd175: sqrt_out <= 22194170;
                10'd176: sqrt_out <= 22257492;
                10'd177: sqrt_out <= 22320634;
                10'd178: sqrt_out <= 22383597;
                10'd179: sqrt_out <= 22446385;
                10'd180: sqrt_out <= 22508997;
                10'd181: sqrt_out <= 22571435;
                10'd182: sqrt_out <= 22633701;
                10'd183: sqrt_out <= 22695797;
                10'd184: sqrt_out <= 22757723;
                10'd185: sqrt_out <= 22819480;
                10'd186: sqrt_out <= 22881072;
                10'd187: sqrt_out <= 22942497;
                10'd188: sqrt_out <= 23003759;
                10'd189: sqrt_out <= 23064858;
                10'd190: sqrt_out <= 23125796;
                10'd191: sqrt_out <= 23186573;
                10'd192: sqrt_out <= 23247192;
                10'd193: sqrt_out <= 23307653;
                10'd194: sqrt_out <= 23367957;
                10'd195: sqrt_out <= 23428107;
                10'd196: sqrt_out <= 23488102;
                10'd197: sqrt_out <= 23547944;
                10'd198: sqrt_out <= 23607635;
                10'd199: sqrt_out <= 23667175;
                10'd200: sqrt_out <= 23726566;
                10'd201: sqrt_out <= 23785808;
                10'd202: sqrt_out <= 23844904;
                10'd203: sqrt_out <= 23903853;
                10'd204: sqrt_out <= 23962657;
                10'd205: sqrt_out <= 24021317;
                10'd206: sqrt_out <= 24079834;
                10'd207: sqrt_out <= 24138210;
                10'd208: sqrt_out <= 24196445;
                10'd209: sqrt_out <= 24254539;
                10'd210: sqrt_out <= 24312495;
                10'd211: sqrt_out <= 24370313;
                10'd212: sqrt_out <= 24427995;
                10'd213: sqrt_out <= 24485540;
                10'd214: sqrt_out <= 24542951;
                10'd215: sqrt_out <= 24600227;
                10'd216: sqrt_out <= 24657371;
                10'd217: sqrt_out <= 24714382;
                10'd218: sqrt_out <= 24771262;
                10'd219: sqrt_out <= 24828012;
                10'd220: sqrt_out <= 24884632;
                10'd221: sqrt_out <= 24941124;
                10'd222: sqrt_out <= 24997488;
                10'd223: sqrt_out <= 25053726;
                10'd224: sqrt_out <= 25109837;
                10'd225: sqrt_out <= 25165824;
                10'd226: sqrt_out <= 25221686;
                10'd227: sqrt_out <= 25277424;
                10'd228: sqrt_out <= 25333040;
                10'd229: sqrt_out <= 25388534;
                10'd230: sqrt_out <= 25443907;
                10'd231: sqrt_out <= 25499160;
                10'd232: sqrt_out <= 25554294;
                10'd233: sqrt_out <= 25609308;
                10'd234: sqrt_out <= 25664205;
                10'd235: sqrt_out <= 25718985;
                10'd236: sqrt_out <= 25773648;
                10'd237: sqrt_out <= 25828195;
                10'd238: sqrt_out <= 25882628;
                10'd239: sqrt_out <= 25936946;
                10'd240: sqrt_out <= 25991151;
                10'd241: sqrt_out <= 26045243;
                10'd242: sqrt_out <= 26099223;
                10'd243: sqrt_out <= 26153091;
                10'd244: sqrt_out <= 26206849;
                10'd245: sqrt_out <= 26260496;
                10'd246: sqrt_out <= 26314035;
                10'd247: sqrt_out <= 26367464;
                10'd248: sqrt_out <= 26420786;
                10'd249: sqrt_out <= 26474000;
                10'd250: sqrt_out <= 26527107;
                10'd251: sqrt_out <= 26580108;
                10'd252: sqrt_out <= 26633004;
                10'd253: sqrt_out <= 26685795;
                10'd254: sqrt_out <= 26738482;
                10'd255: sqrt_out <= 26791065;
                10'd256: sqrt_out <= 26843545;
                10'd257: sqrt_out <= 26895923;
                10'd258: sqrt_out <= 26948199;
                10'd259: sqrt_out <= 27000373;
                10'd260: sqrt_out <= 27052447;
                10'd261: sqrt_out <= 27104421;
                10'd262: sqrt_out <= 27156296;
                10'd263: sqrt_out <= 27208072;
                10'd264: sqrt_out <= 27259749;
                10'd265: sqrt_out <= 27311328;
                10'd266: sqrt_out <= 27362811;
                10'd267: sqrt_out <= 27414196;
                10'd268: sqrt_out <= 27465486;
                10'd269: sqrt_out <= 27516680;
                10'd270: sqrt_out <= 27567778;
                10'd271: sqrt_out <= 27618783;
                10'd272: sqrt_out <= 27669693;
                10'd273: sqrt_out <= 27720510;
                10'd274: sqrt_out <= 27771233;
                10'd275: sqrt_out <= 27821865;
                10'd276: sqrt_out <= 27872404;
                10'd277: sqrt_out <= 27922852;
                10'd278: sqrt_out <= 27973209;
                10'd279: sqrt_out <= 28023475;
                10'd280: sqrt_out <= 28073651;
                10'd281: sqrt_out <= 28123738;
                10'd282: sqrt_out <= 28173736;
                10'd283: sqrt_out <= 28223645;
                10'd284: sqrt_out <= 28273466;
                10'd285: sqrt_out <= 28323200;
                10'd286: sqrt_out <= 28372846;
                10'd287: sqrt_out <= 28422406;
                10'd288: sqrt_out <= 28471879;
                10'd289: sqrt_out <= 28521267;
                10'd290: sqrt_out <= 28570569;
                10'd291: sqrt_out <= 28619786;
                10'd292: sqrt_out <= 28668919;
                10'd293: sqrt_out <= 28717967;
                10'd294: sqrt_out <= 28766932;
                10'd295: sqrt_out <= 28815814;
                10'd296: sqrt_out <= 28864613;
                10'd297: sqrt_out <= 28913330;
                10'd298: sqrt_out <= 28961965;
                10'd299: sqrt_out <= 29010518;
                10'd300: sqrt_out <= 29058990;
                10'd301: sqrt_out <= 29107381;
                10'd302: sqrt_out <= 29155692;
                10'd303: sqrt_out <= 29203924;
                10'd304: sqrt_out <= 29252075;
                10'd305: sqrt_out <= 29300148;
                10'd306: sqrt_out <= 29348141;
                10'd307: sqrt_out <= 29396057;
                10'd308: sqrt_out <= 29443894;
                10'd309: sqrt_out <= 29491654;
                10'd310: sqrt_out <= 29539336;
                10'd311: sqrt_out <= 29586942;
                10'd312: sqrt_out <= 29634471;
                10'd313: sqrt_out <= 29681925;
                10'd314: sqrt_out <= 29729302;
                10'd315: sqrt_out <= 29776604;
                10'd316: sqrt_out <= 29823831;
                10'd317: sqrt_out <= 29870983;
                10'd318: sqrt_out <= 29918061;
                10'd319: sqrt_out <= 29965065;
                10'd320: sqrt_out <= 30011996;
                10'd321: sqrt_out <= 30058853;
                10'd322: sqrt_out <= 30105637;
                10'd323: sqrt_out <= 30152349;
                10'd324: sqrt_out <= 30198988;
                10'd325: sqrt_out <= 30245556;
                10'd326: sqrt_out <= 30292052;
                10'd327: sqrt_out <= 30338476;
                10'd328: sqrt_out <= 30384830;
                10'd329: sqrt_out <= 30431113;
                10'd330: sqrt_out <= 30477326;
                10'd331: sqrt_out <= 30523469;
                10'd332: sqrt_out <= 30569542;
                10'd333: sqrt_out <= 30615546;
                10'd334: sqrt_out <= 30661481;
                10'd335: sqrt_out <= 30707347;
                10'd336: sqrt_out <= 30753144;
                10'd337: sqrt_out <= 30798874;
                10'd338: sqrt_out <= 30844536;
                10'd339: sqrt_out <= 30890130;
                10'd340: sqrt_out <= 30935657;
                10'd341: sqrt_out <= 30981117;
                10'd342: sqrt_out <= 31026511;
                10'd343: sqrt_out <= 31071838;
                10'd344: sqrt_out <= 31117100;
                10'd345: sqrt_out <= 31162295;
                10'd346: sqrt_out <= 31207425;
                10'd347: sqrt_out <= 31252490;
                10'd348: sqrt_out <= 31297490;
                10'd349: sqrt_out <= 31342426;
                10'd350: sqrt_out <= 31387297;
                10'd351: sqrt_out <= 31432104;
                10'd352: sqrt_out <= 31476847;
                10'd353: sqrt_out <= 31521527;
                10'd354: sqrt_out <= 31566143;
                10'd355: sqrt_out <= 31610697;
                10'd356: sqrt_out <= 31655187;
                10'd357: sqrt_out <= 31699616;
                10'd358: sqrt_out <= 31743982;
                10'd359: sqrt_out <= 31788286;
                10'd360: sqrt_out <= 31832529;
                10'd361: sqrt_out <= 31876710;
                10'd362: sqrt_out <= 31920830;
                10'd363: sqrt_out <= 31964889;
                10'd364: sqrt_out <= 32008888;
                10'd365: sqrt_out <= 32052826;
                10'd366: sqrt_out <= 32096704;
                10'd367: sqrt_out <= 32140522;
                10'd368: sqrt_out <= 32184280;
                10'd369: sqrt_out <= 32227979;
                10'd370: sqrt_out <= 32271619;
                10'd371: sqrt_out <= 32315200;
                10'd372: sqrt_out <= 32358722;
                10'd373: sqrt_out <= 32402186;
                10'd374: sqrt_out <= 32445591;
                10'd375: sqrt_out <= 32488939;
                10'd376: sqrt_out <= 32532228;
                10'd377: sqrt_out <= 32575461;
                10'd378: sqrt_out <= 32618635;
                10'd379: sqrt_out <= 32661753;
                10'd380: sqrt_out <= 32704814;
                10'd381: sqrt_out <= 32747819;
                10'd382: sqrt_out <= 32790767;
                10'd383: sqrt_out <= 32833658;
                10'd384: sqrt_out <= 32876494;
                10'd385: sqrt_out <= 32919274;
                10'd386: sqrt_out <= 32961999;
                10'd387: sqrt_out <= 33004668;
                10'd388: sqrt_out <= 33047282;
                10'd389: sqrt_out <= 33089842;
                10'd390: sqrt_out <= 33132346;
                10'd391: sqrt_out <= 33174797;
                10'd392: sqrt_out <= 33217192;
                10'd393: sqrt_out <= 33259534;
                10'd394: sqrt_out <= 33301822;
                10'd395: sqrt_out <= 33344057;
                10'd396: sqrt_out <= 33386238;
                10'd397: sqrt_out <= 33428366;
                10'd398: sqrt_out <= 33470440;
                10'd399: sqrt_out <= 33512462;
                10'd400: sqrt_out <= 33554432;
                10'd401: sqrt_out <= 33596348;
                10'd402: sqrt_out <= 33638213;
                10'd403: sqrt_out <= 33680026;
                10'd404: sqrt_out <= 33721786;
                10'd405: sqrt_out <= 33763495;
                10'd406: sqrt_out <= 33805153;
                10'd407: sqrt_out <= 33846759;
                10'd408: sqrt_out <= 33888315;
                10'd409: sqrt_out <= 33929819;
                10'd410: sqrt_out <= 33971273;
                10'd411: sqrt_out <= 34012676;
                10'd412: sqrt_out <= 34054029;
                10'd413: sqrt_out <= 34095331;
                10'd414: sqrt_out <= 34136584;
                10'd415: sqrt_out <= 34177787;
                10'd416: sqrt_out <= 34218940;
                10'd417: sqrt_out <= 34260044;
                10'd418: sqrt_out <= 34301099;
                10'd419: sqrt_out <= 34342104;
                10'd420: sqrt_out <= 34383061;
                10'd421: sqrt_out <= 34423969;
                10'd422: sqrt_out <= 34464828;
                10'd423: sqrt_out <= 34505639;
                10'd424: sqrt_out <= 34546402;
                10'd425: sqrt_out <= 34587116;
                10'd426: sqrt_out <= 34627783;
                10'd427: sqrt_out <= 34668402;
                10'd428: sqrt_out <= 34708974;
                10'd429: sqrt_out <= 34749498;
                10'd430: sqrt_out <= 34789975;
                10'd431: sqrt_out <= 34830405;
                10'd432: sqrt_out <= 34870788;
                10'd433: sqrt_out <= 34911125;
                10'd434: sqrt_out <= 34951414;
                10'd435: sqrt_out <= 34991658;
                10'd436: sqrt_out <= 35031855;
                10'd437: sqrt_out <= 35072006;
                10'd438: sqrt_out <= 35112111;
                10'd439: sqrt_out <= 35152171;
                10'd440: sqrt_out <= 35192185;
                10'd441: sqrt_out <= 35232153;
                10'd442: sqrt_out <= 35272076;
                10'd443: sqrt_out <= 35311954;
                10'd444: sqrt_out <= 35351787;
                10'd445: sqrt_out <= 35391575;
                10'd446: sqrt_out <= 35431319;
                10'd447: sqrt_out <= 35471018;
                10'd448: sqrt_out <= 35510672;
                10'd449: sqrt_out <= 35550283;
                10'd450: sqrt_out <= 35589849;
                10'd451: sqrt_out <= 35629371;
                10'd452: sqrt_out <= 35668850;
                10'd453: sqrt_out <= 35708285;
                10'd454: sqrt_out <= 35747676;
                10'd455: sqrt_out <= 35787024;
                10'd456: sqrt_out <= 35826329;
                10'd457: sqrt_out <= 35865591;
                10'd458: sqrt_out <= 35904810;
                10'd459: sqrt_out <= 35943986;
                10'd460: sqrt_out <= 35983119;
                10'd461: sqrt_out <= 36022210;
                10'd462: sqrt_out <= 36061258;
                10'd463: sqrt_out <= 36100265;
                10'd464: sqrt_out <= 36139229;
                10'd465: sqrt_out <= 36178151;
                10'd466: sqrt_out <= 36217031;
                10'd467: sqrt_out <= 36255870;
                10'd468: sqrt_out <= 36294667;
                10'd469: sqrt_out <= 36333423;
                10'd470: sqrt_out <= 36372137;
                10'd471: sqrt_out <= 36410810;
                10'd472: sqrt_out <= 36449442;
                10'd473: sqrt_out <= 36488034;
                10'd474: sqrt_out <= 36526584;
                10'd475: sqrt_out <= 36565094;
                10'd476: sqrt_out <= 36603563;
                10'd477: sqrt_out <= 36641992;
                10'd478: sqrt_out <= 36680381;
                10'd479: sqrt_out <= 36718730;
                10'd480: sqrt_out <= 36757038;
                10'd481: sqrt_out <= 36795307;
                10'd482: sqrt_out <= 36833536;
                10'd483: sqrt_out <= 36871725;
                10'd484: sqrt_out <= 36909875;
                10'd485: sqrt_out <= 36947985;
                10'd486: sqrt_out <= 36986056;
                10'd487: sqrt_out <= 37024088;
                10'd488: sqrt_out <= 37062081;
                10'd489: sqrt_out <= 37100035;
                10'd490: sqrt_out <= 37137950;
                10'd491: sqrt_out <= 37175827;
                10'd492: sqrt_out <= 37213665;
                10'd493: sqrt_out <= 37251464;
                10'd494: sqrt_out <= 37289226;
                10'd495: sqrt_out <= 37326949;
                10'd496: sqrt_out <= 37364634;
                10'd497: sqrt_out <= 37402281;
                10'd498: sqrt_out <= 37439890;
                10'd499: sqrt_out <= 37477461;
                10'd500: sqrt_out <= 37514995;
                10'd501: sqrt_out <= 37552491;
                10'd502: sqrt_out <= 37589950;
                10'd503: sqrt_out <= 37627372;
                10'd504: sqrt_out <= 37664756;
                10'd505: sqrt_out <= 37702103;
                10'd506: sqrt_out <= 37739414;
                10'd507: sqrt_out <= 37776687;
                10'd508: sqrt_out <= 37813924;
                10'd509: sqrt_out <= 37851124;
                10'd510: sqrt_out <= 37888288;
                10'd511: sqrt_out <= 37925415;
                10'd512: sqrt_out <= 37962506;
                10'd513: sqrt_out <= 37999560;
                10'd514: sqrt_out <= 38036579;
                10'd515: sqrt_out <= 38073562;
                10'd516: sqrt_out <= 38110508;
                10'd517: sqrt_out <= 38147419;
                10'd518: sqrt_out <= 38184294;
                10'd519: sqrt_out <= 38221134;
                10'd520: sqrt_out <= 38257938;
                10'd521: sqrt_out <= 38294707;
                10'd522: sqrt_out <= 38331441;
                10'd523: sqrt_out <= 38368139;
                10'd524: sqrt_out <= 38404802;
                10'd525: sqrt_out <= 38441431;
                10'd526: sqrt_out <= 38478024;
                10'd527: sqrt_out <= 38514583;
                10'd528: sqrt_out <= 38551107;
                10'd529: sqrt_out <= 38587596;
                10'd530: sqrt_out <= 38624051;
                10'd531: sqrt_out <= 38660472;
                10'd532: sqrt_out <= 38696858;
                10'd533: sqrt_out <= 38733210;
                10'd534: sqrt_out <= 38769528;
                10'd535: sqrt_out <= 38805813;
                10'd536: sqrt_out <= 38842063;
                10'd537: sqrt_out <= 38878279;
                10'd538: sqrt_out <= 38914462;
                10'd539: sqrt_out <= 38950611;
                10'd540: sqrt_out <= 38986726;
                10'd541: sqrt_out <= 39022809;
                10'd542: sqrt_out <= 39058857;
                10'd543: sqrt_out <= 39094873;
                10'd544: sqrt_out <= 39130855;
                10'd545: sqrt_out <= 39166805;
                10'd546: sqrt_out <= 39202721;
                10'd547: sqrt_out <= 39238605;
                10'd548: sqrt_out <= 39274455;
                10'd549: sqrt_out <= 39310273;
                10'd550: sqrt_out <= 39346059;
                10'd551: sqrt_out <= 39381812;
                10'd552: sqrt_out <= 39417532;
                10'd553: sqrt_out <= 39453220;
                10'd554: sqrt_out <= 39488876;
                10'd555: sqrt_out <= 39524500;
                10'd556: sqrt_out <= 39560091;
                10'd557: sqrt_out <= 39595651;
                10'd558: sqrt_out <= 39631179;
                10'd559: sqrt_out <= 39666675;
                10'd560: sqrt_out <= 39702139;
                10'd561: sqrt_out <= 39737571;
                10'd562: sqrt_out <= 39772972;
                10'd563: sqrt_out <= 39808342;
                10'd564: sqrt_out <= 39843680;
                10'd565: sqrt_out <= 39878987;
                10'd566: sqrt_out <= 39914262;
                10'd567: sqrt_out <= 39949507;
                10'd568: sqrt_out <= 39984720;
                10'd569: sqrt_out <= 40019902;
                10'd570: sqrt_out <= 40055054;
                10'd571: sqrt_out <= 40090174;
                10'd572: sqrt_out <= 40125264;
                10'd573: sqrt_out <= 40160323;
                10'd574: sqrt_out <= 40195352;
                10'd575: sqrt_out <= 40230350;
                10'd576: sqrt_out <= 40265318;
                10'd577: sqrt_out <= 40300255;
                10'd578: sqrt_out <= 40335162;
                10'd579: sqrt_out <= 40370039;
                10'd580: sqrt_out <= 40404886;
                10'd581: sqrt_out <= 40439703;
                10'd582: sqrt_out <= 40474490;
                10'd583: sqrt_out <= 40509247;
                10'd584: sqrt_out <= 40543974;
                10'd585: sqrt_out <= 40578671;
                10'd586: sqrt_out <= 40613339;
                10'd587: sqrt_out <= 40647977;
                10'd588: sqrt_out <= 40682586;
                10'd589: sqrt_out <= 40717166;
                10'd590: sqrt_out <= 40751716;
                10'd591: sqrt_out <= 40786236;
                10'd592: sqrt_out <= 40820728;
                10'd593: sqrt_out <= 40855190;
                10'd594: sqrt_out <= 40889624;
                10'd595: sqrt_out <= 40924028;
                10'd596: sqrt_out <= 40958404;
                10'd597: sqrt_out <= 40992750;
                10'd598: sqrt_out <= 41027068;
                10'd599: sqrt_out <= 41061357;
                10'd600: sqrt_out <= 41095618;
                10'd601: sqrt_out <= 41129850;
                10'd602: sqrt_out <= 41164054;
                10'd603: sqrt_out <= 41198229;
                10'd604: sqrt_out <= 41232376;
                10'd605: sqrt_out <= 41266494;
                10'd606: sqrt_out <= 41300585;
                10'd607: sqrt_out <= 41334647;
                10'd608: sqrt_out <= 41368682;
                10'd609: sqrt_out <= 41402688;
                10'd610: sqrt_out <= 41436666;
                10'd611: sqrt_out <= 41470617;
                10'd612: sqrt_out <= 41504540;
                10'd613: sqrt_out <= 41538435;
                10'd614: sqrt_out <= 41572302;
                10'd615: sqrt_out <= 41606142;
                10'd616: sqrt_out <= 41639955;
                10'd617: sqrt_out <= 41673740;
                10'd618: sqrt_out <= 41707497;
                10'd619: sqrt_out <= 41741227;
                10'd620: sqrt_out <= 41774930;
                10'd621: sqrt_out <= 41808606;
                10'd622: sqrt_out <= 41842255;
                10'd623: sqrt_out <= 41875877;
                10'd624: sqrt_out <= 41909472;
                10'd625: sqrt_out <= 41943040;
                10'd626: sqrt_out <= 41976581;
                10'd627: sqrt_out <= 42010095;
                10'd628: sqrt_out <= 42043582;
                10'd629: sqrt_out <= 42077043;
                10'd630: sqrt_out <= 42110477;
                10'd631: sqrt_out <= 42143885;
                10'd632: sqrt_out <= 42177267;
                10'd633: sqrt_out <= 42210621;
                10'd634: sqrt_out <= 42243950;
                10'd635: sqrt_out <= 42277252;
                10'd636: sqrt_out <= 42310528;
                10'd637: sqrt_out <= 42343778;
                10'd638: sqrt_out <= 42377002;
                10'd639: sqrt_out <= 42410200;
                10'd640: sqrt_out <= 42443372;
                10'd641: sqrt_out <= 42476518;
                10'd642: sqrt_out <= 42509638;
                10'd643: sqrt_out <= 42542732;
                10'd644: sqrt_out <= 42575801;
                10'd645: sqrt_out <= 42608844;
                10'd646: sqrt_out <= 42641861;
                10'd647: sqrt_out <= 42674853;
                10'd648: sqrt_out <= 42707819;
                10'd649: sqrt_out <= 42740760;
                10'd650: sqrt_out <= 42773675;
                10'd651: sqrt_out <= 42806566;
                10'd652: sqrt_out <= 42839430;
                10'd653: sqrt_out <= 42872270;
                10'd654: sqrt_out <= 42905085;
                10'd655: sqrt_out <= 42937874;
                10'd656: sqrt_out <= 42970639;
                10'd657: sqrt_out <= 43003378;
                10'd658: sqrt_out <= 43036093;
                10'd659: sqrt_out <= 43068783;
                10'd660: sqrt_out <= 43101448;
                10'd661: sqrt_out <= 43134088;
                10'd662: sqrt_out <= 43166704;
                10'd663: sqrt_out <= 43199295;
                10'd664: sqrt_out <= 43231861;
                10'd665: sqrt_out <= 43264403;
                10'd666: sqrt_out <= 43296920;
                10'd667: sqrt_out <= 43329413;
                10'd668: sqrt_out <= 43361882;
                10'd669: sqrt_out <= 43394326;
                10'd670: sqrt_out <= 43426746;
                10'd671: sqrt_out <= 43459142;
                10'd672: sqrt_out <= 43491514;
                10'd673: sqrt_out <= 43523862;
                10'd674: sqrt_out <= 43556186;
                10'd675: sqrt_out <= 43588485;
                10'd676: sqrt_out <= 43620761;
                10'd677: sqrt_out <= 43653013;
                10'd678: sqrt_out <= 43685241;
                10'd679: sqrt_out <= 43717446;
                10'd680: sqrt_out <= 43749626;
                10'd681: sqrt_out <= 43781783;
                10'd682: sqrt_out <= 43813917;
                10'd683: sqrt_out <= 43846027;
                10'd684: sqrt_out <= 43878113;
                10'd685: sqrt_out <= 43910176;
                10'd686: sqrt_out <= 43942215;
                10'd687: sqrt_out <= 43974232;
                10'd688: sqrt_out <= 44006225;
                10'd689: sqrt_out <= 44038194;
                10'd690: sqrt_out <= 44070141;
                10'd691: sqrt_out <= 44102064;
                10'd692: sqrt_out <= 44133964;
                10'd693: sqrt_out <= 44165841;
                10'd694: sqrt_out <= 44197696;
                10'd695: sqrt_out <= 44229527;
                10'd696: sqrt_out <= 44261335;
                10'd697: sqrt_out <= 44293121;
                10'd698: sqrt_out <= 44324883;
                10'd699: sqrt_out <= 44356623;
                10'd700: sqrt_out <= 44388341;
                10'd701: sqrt_out <= 44420035;
                10'd702: sqrt_out <= 44451707;
                10'd703: sqrt_out <= 44483357;
                10'd704: sqrt_out <= 44514984;
                10'd705: sqrt_out <= 44546588;
                10'd706: sqrt_out <= 44578171;
                10'd707: sqrt_out <= 44609730;
                10'd708: sqrt_out <= 44641268;
                10'd709: sqrt_out <= 44672783;
                10'd710: sqrt_out <= 44704276;
                10'd711: sqrt_out <= 44735747;
                10'd712: sqrt_out <= 44767195;
                10'd713: sqrt_out <= 44798622;
                10'd714: sqrt_out <= 44830027;
                10'd715: sqrt_out <= 44861409;
                10'd716: sqrt_out <= 44892770;
                10'd717: sqrt_out <= 44924109;
                10'd718: sqrt_out <= 44955426;
                10'd719: sqrt_out <= 44986721;
                10'd720: sqrt_out <= 45017994;
                10'd721: sqrt_out <= 45049246;
                10'd722: sqrt_out <= 45080476;
                10'd723: sqrt_out <= 45111684;
                10'd724: sqrt_out <= 45142871;
                10'd725: sqrt_out <= 45174036;
                10'd726: sqrt_out <= 45205180;
                10'd727: sqrt_out <= 45236302;
                10'd728: sqrt_out <= 45267403;
                10'd729: sqrt_out <= 45298483;
                10'd730: sqrt_out <= 45329541;
                10'd731: sqrt_out <= 45360578;
                10'd732: sqrt_out <= 45391594;
                10'd733: sqrt_out <= 45422588;
                10'd734: sqrt_out <= 45453562;
                10'd735: sqrt_out <= 45484514;
                10'd736: sqrt_out <= 45515446;
                10'd737: sqrt_out <= 45546356;
                10'd738: sqrt_out <= 45577245;
                10'd739: sqrt_out <= 45608114;
                10'd740: sqrt_out <= 45638961;
                10'd741: sqrt_out <= 45669788;
                10'd742: sqrt_out <= 45700594;
                10'd743: sqrt_out <= 45731379;
                10'd744: sqrt_out <= 45762144;
                10'd745: sqrt_out <= 45792887;
                10'd746: sqrt_out <= 45823611;
                10'd747: sqrt_out <= 45854313;
                10'd748: sqrt_out <= 45884995;
                10'd749: sqrt_out <= 45915657;
                10'd750: sqrt_out <= 45946298;
                10'd751: sqrt_out <= 45976918;
                10'd752: sqrt_out <= 46007519;
                10'd753: sqrt_out <= 46038099;
                10'd754: sqrt_out <= 46068658;
                10'd755: sqrt_out <= 46099198;
                10'd756: sqrt_out <= 46129717;
                10'd757: sqrt_out <= 46160216;
                10'd758: sqrt_out <= 46190695;
                10'd759: sqrt_out <= 46221153;
                10'd760: sqrt_out <= 46251592;
                10'd761: sqrt_out <= 46282011;
                10'd762: sqrt_out <= 46312410;
                10'd763: sqrt_out <= 46342788;
                10'd764: sqrt_out <= 46373147;
                10'd765: sqrt_out <= 46403486;
                10'd766: sqrt_out <= 46433805;
                10'd767: sqrt_out <= 46464105;
                10'd768: sqrt_out <= 46494384;
                10'd769: sqrt_out <= 46524644;
                10'd770: sqrt_out <= 46554885;
                10'd771: sqrt_out <= 46585105;
                10'd772: sqrt_out <= 46615306;
                10'd773: sqrt_out <= 46645488;
                10'd774: sqrt_out <= 46675650;
                10'd775: sqrt_out <= 46705792;
                10'd776: sqrt_out <= 46735915;
                10'd777: sqrt_out <= 46766019;
                10'd778: sqrt_out <= 46796103;
                10'd779: sqrt_out <= 46826168;
                10'd780: sqrt_out <= 46856214;
                10'd781: sqrt_out <= 46886240;
                10'd782: sqrt_out <= 46916247;
                10'd783: sqrt_out <= 46946235;
                10'd784: sqrt_out <= 46976204;
                10'd785: sqrt_out <= 47006154;
                10'd786: sqrt_out <= 47036085;
                10'd787: sqrt_out <= 47065996;
                10'd788: sqrt_out <= 47095889;
                10'd789: sqrt_out <= 47125763;
                10'd790: sqrt_out <= 47155618;
                10'd791: sqrt_out <= 47185453;
                10'd792: sqrt_out <= 47215270;
                10'd793: sqrt_out <= 47245069;
                10'd794: sqrt_out <= 47274848;
                10'd795: sqrt_out <= 47304609;
                10'd796: sqrt_out <= 47334351;
                10'd797: sqrt_out <= 47364074;
                10'd798: sqrt_out <= 47393779;
                10'd799: sqrt_out <= 47423465;
                10'd800: sqrt_out <= 47453132;
                10'd801: sqrt_out <= 47482781;
                10'd802: sqrt_out <= 47512412;
                10'd803: sqrt_out <= 47542024;
                10'd804: sqrt_out <= 47571617;
                10'd805: sqrt_out <= 47601192;
                10'd806: sqrt_out <= 47630749;
                10'd807: sqrt_out <= 47660288;
                10'd808: sqrt_out <= 47689808;
                10'd809: sqrt_out <= 47719310;
                10'd810: sqrt_out <= 47748793;
                10'd811: sqrt_out <= 47778259;
                10'd812: sqrt_out <= 47807706;
                10'd813: sqrt_out <= 47837135;
                10'd814: sqrt_out <= 47866546;
                10'd815: sqrt_out <= 47895939;
                10'd816: sqrt_out <= 47925314;
                10'd817: sqrt_out <= 47954671;
                10'd818: sqrt_out <= 47984010;
                10'd819: sqrt_out <= 48013332;
                10'd820: sqrt_out <= 48042635;
                10'd821: sqrt_out <= 48071920;
                10'd822: sqrt_out <= 48101188;
                10'd823: sqrt_out <= 48130437;
                10'd824: sqrt_out <= 48159669;
                10'd825: sqrt_out <= 48188884;
                10'd826: sqrt_out <= 48218080;
                10'd827: sqrt_out <= 48247259;
                10'd828: sqrt_out <= 48276420;
                10'd829: sqrt_out <= 48305564;
                10'd830: sqrt_out <= 48334690;
                10'd831: sqrt_out <= 48363799;
                10'd832: sqrt_out <= 48392890;
                10'd833: sqrt_out <= 48421963;
                10'd834: sqrt_out <= 48451019;
                10'd835: sqrt_out <= 48480058;
                10'd836: sqrt_out <= 48509079;
                10'd837: sqrt_out <= 48538083;
                10'd838: sqrt_out <= 48567070;
                10'd839: sqrt_out <= 48596039;
                10'd840: sqrt_out <= 48624991;
                10'd841: sqrt_out <= 48653926;
                10'd842: sqrt_out <= 48682844;
                10'd843: sqrt_out <= 48711744;
                10'd844: sqrt_out <= 48740627;
                10'd845: sqrt_out <= 48769494;
                10'd846: sqrt_out <= 48798343;
                10'd847: sqrt_out <= 48827175;
                10'd848: sqrt_out <= 48855990;
                10'd849: sqrt_out <= 48884788;
                10'd850: sqrt_out <= 48913569;
                10'd851: sqrt_out <= 48942333;
                10'd852: sqrt_out <= 48971081;
                10'd853: sqrt_out <= 48999811;
                10'd854: sqrt_out <= 49028525;
                10'd855: sqrt_out <= 49057222;
                10'd856: sqrt_out <= 49085902;
                10'd857: sqrt_out <= 49114565;
                10'd858: sqrt_out <= 49143212;
                10'd859: sqrt_out <= 49171842;
                10'd860: sqrt_out <= 49200455;
                10'd861: sqrt_out <= 49229051;
                10'd862: sqrt_out <= 49257631;
                10'd863: sqrt_out <= 49286195;
                10'd864: sqrt_out <= 49314742;
                10'd865: sqrt_out <= 49343272;
                10'd866: sqrt_out <= 49371786;
                10'd867: sqrt_out <= 49400283;
                10'd868: sqrt_out <= 49428764;
                10'd869: sqrt_out <= 49457229;
                10'd870: sqrt_out <= 49485677;
                10'd871: sqrt_out <= 49514109;
                10'd872: sqrt_out <= 49542525;
                10'd873: sqrt_out <= 49570924;
                10'd874: sqrt_out <= 49599307;
                10'd875: sqrt_out <= 49627674;
                10'd876: sqrt_out <= 49656024;
                10'd877: sqrt_out <= 49684359;
                10'd878: sqrt_out <= 49712677;
                10'd879: sqrt_out <= 49740979;
                10'd880: sqrt_out <= 49769265;
                10'd881: sqrt_out <= 49797535;
                10'd882: sqrt_out <= 49825789;
                10'd883: sqrt_out <= 49854027;
                10'd884: sqrt_out <= 49882249;
                10'd885: sqrt_out <= 49910455;
                10'd886: sqrt_out <= 49938645;
                10'd887: sqrt_out <= 49966819;
                10'd888: sqrt_out <= 49994977;
                10'd889: sqrt_out <= 50023120;
                10'd890: sqrt_out <= 50051246;
                10'd891: sqrt_out <= 50079357;
                10'd892: sqrt_out <= 50107452;
                10'd893: sqrt_out <= 50135531;
                10'd894: sqrt_out <= 50163595;
                10'd895: sqrt_out <= 50191643;
                10'd896: sqrt_out <= 50219675;
                10'd897: sqrt_out <= 50247691;
                10'd898: sqrt_out <= 50275692;
                10'd899: sqrt_out <= 50303678;
                10'd900: sqrt_out <= 50331648;
                10'd901: sqrt_out <= 50359602;
                10'd902: sqrt_out <= 50387541;
                10'd903: sqrt_out <= 50415464;
                10'd904: sqrt_out <= 50443372;
                10'd905: sqrt_out <= 50471264;
                10'd906: sqrt_out <= 50499141;
                10'd907: sqrt_out <= 50527003;
                10'd908: sqrt_out <= 50554849;
                10'd909: sqrt_out <= 50582680;
                10'd910: sqrt_out <= 50610495;
                10'd911: sqrt_out <= 50638296;
                10'd912: sqrt_out <= 50666081;
                10'd913: sqrt_out <= 50693851;
                10'd914: sqrt_out <= 50721605;
                10'd915: sqrt_out <= 50749345;
                10'd916: sqrt_out <= 50777069;
                10'd917: sqrt_out <= 50804778;
                10'd918: sqrt_out <= 50832472;
                10'd919: sqrt_out <= 50860151;
                10'd920: sqrt_out <= 50887815;
                10'd921: sqrt_out <= 50915464;
                10'd922: sqrt_out <= 50943098;
                10'd923: sqrt_out <= 50970717;
                10'd924: sqrt_out <= 50998321;
                10'd925: sqrt_out <= 51025910;
                10'd926: sqrt_out <= 51053484;
                10'd927: sqrt_out <= 51081043;
                10'd928: sqrt_out <= 51108588;
                10'd929: sqrt_out <= 51136117;
                10'd930: sqrt_out <= 51163632;
                10'd931: sqrt_out <= 51191132;
                10'd932: sqrt_out <= 51218617;
                10'd933: sqrt_out <= 51246087;
                10'd934: sqrt_out <= 51273543;
                10'd935: sqrt_out <= 51300984;
                10'd936: sqrt_out <= 51328411;
                10'd937: sqrt_out <= 51355822;
                10'd938: sqrt_out <= 51383219;
                10'd939: sqrt_out <= 51410602;
                10'd940: sqrt_out <= 51437970;
                10'd941: sqrt_out <= 51465323;
                10'd942: sqrt_out <= 51492662;
                10'd943: sqrt_out <= 51519986;
                10'd944: sqrt_out <= 51547296;
                10'd945: sqrt_out <= 51574591;
                10'd946: sqrt_out <= 51601872;
                10'd947: sqrt_out <= 51629139;
                10'd948: sqrt_out <= 51656391;
                10'd949: sqrt_out <= 51683629;
                10'd950: sqrt_out <= 51710852;
                10'd951: sqrt_out <= 51738061;
                10'd952: sqrt_out <= 51765256;
                10'd953: sqrt_out <= 51792436;
                10'd954: sqrt_out <= 51819603;
                10'd955: sqrt_out <= 51846755;
                10'd956: sqrt_out <= 51873893;
                10'd957: sqrt_out <= 51901016;
                10'd958: sqrt_out <= 51928126;
                10'd959: sqrt_out <= 51955221;
                10'd960: sqrt_out <= 51982302;
                10'd961: sqrt_out <= 52009369;
                10'd962: sqrt_out <= 52036422;
                10'd963: sqrt_out <= 52063461;
                10'd964: sqrt_out <= 52090486;
                10'd965: sqrt_out <= 52117497;
                10'd966: sqrt_out <= 52144494;
                10'd967: sqrt_out <= 52171477;
                10'd968: sqrt_out <= 52198446;
                10'd969: sqrt_out <= 52225401;
                10'd970: sqrt_out <= 52252342;
                10'd971: sqrt_out <= 52279269;
                10'd972: sqrt_out <= 52306182;
                10'd973: sqrt_out <= 52333082;
                10'd974: sqrt_out <= 52359968;
                10'd975: sqrt_out <= 52386840;
                10'd976: sqrt_out <= 52413698;
                10'd977: sqrt_out <= 52440542;
                10'd978: sqrt_out <= 52467373;
                10'd979: sqrt_out <= 52494190;
                10'd980: sqrt_out <= 52520993;
                10'd981: sqrt_out <= 52547783;
                10'd982: sqrt_out <= 52574559;
                10'd983: sqrt_out <= 52601321;
                10'd984: sqrt_out <= 52628070;
                10'd985: sqrt_out <= 52654805;
                10'd986: sqrt_out <= 52681526;
                10'd987: sqrt_out <= 52708234;
                10'd988: sqrt_out <= 52734929;
                10'd989: sqrt_out <= 52761610;
                10'd990: sqrt_out <= 52788277;
                10'd991: sqrt_out <= 52814931;
                10'd992: sqrt_out <= 52841572;
                10'd993: sqrt_out <= 52868199;
                10'd994: sqrt_out <= 52894813;
                10'd995: sqrt_out <= 52921413;
                10'd996: sqrt_out <= 52948000;
                10'd997: sqrt_out <= 52974574;
                10'd998: sqrt_out <= 53001134;
                10'd999: sqrt_out <= 53027681;
                10'd1000: sqrt_out <= 53054215;
                default: cos_out <= -32'hFFFFFFFF;
            endcase
        end
    end
endmodule